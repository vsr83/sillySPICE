SIMPLE CIRCUIT WITH VOLTAGE-CONTROLLED VOLTAGE SOURCE
V1 1 0 1
R1 2 1 1
R2 0 2 2
E1 2 0 1 2 3
*FOOOBAR
.dc v1 1 1 2
.end