SIMPLE CIRCUIT WITH VOLTAGE-CONTROLLED CURRENT SOURCE
V1 1 0 1
R1 2 1 1
R2 0 2 1
G1 2 0 1 2 1
*FOOOBAR
.dc v1 1 1 2
.end