SIMPLE CIRCUIT WITH A CURRENT SOURCE
R1   1 0 1
R2   1 0 1
IDC 1 0 1
*FOOOBAR
.dc IDC 0 1 2
.end