SIMPLE CIRCUIT WITH A CURRENT SOURCE
VDC 1 0 1
R1   2 1 1000
C1   0 2 1
*FOOOBAR
.tran 0 1
.end
