SIMPLE CIRCUIT
R1 2 1 1  ; vittumainen vastus
R2 3 2 1
R3 4 3 1
R4 0 4 1
VDC 1 0 4 
*FOOOBAR
.dc VDC 0 1 2
.end