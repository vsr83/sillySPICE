SIMPLE CAPACITIVE CIRCUIT
* Analytical solution can be easily obtained as:

IAC 1 0 PULSE (0 1 0.0001 0.0001 0.0001 0.05 0.1) 
R1   2 1 100
L1   0 2 1

.tran 0 1
.end
