SIMPLE CIRCUIT
R1   2 1 1
VDC  1 0 1
R2   0 2 2
F1   2 0 vdc 3
*FOOOBAR
.dc vdc 0 1 2
.end